ta en pil .
ta ett block .
ta en kon .
ta en blå kon .
ta en röd kon .
ta en blå pil .
ta en röd pil .
hämta ett block .
ta blocket .
ta inte blocket .
ta pilen .
ställ en kon på mitt block .
ställ en kon på hans block .
ställ en kon på hennes block .
ställ en kon på blocket .
hon tar blocket .
hon tar pyramiden .
ställ en blå pil på en blå cirkel .
ställ en röd pil på en blå cirkel .
ställ en lila pil på en blå cirkel .
jag tar ett blått block .
jag tar ett rött block .
ställ blocket på cirkeln .
ställ konen på cirkeln .
ställ pilen på cirkeln .
han ställer det röda blocket på den blåa cirkeln .
han ställer det röda blocket på den röda cirkeln .
han ställer det blå blocket på den röda cirkeln .
han ställer en pil på min cirkel .
han ställer en pil på sin cirkel .
han ställer en pil på hans cirkel .
han ställer en pil på hennes cirkel .
hon ställer sitt block på min blåa cirkel .
hon ställer sitt block på min röda cirkel .
jag ställer konen på cirkeln på hennes blåa cirkel .
jag ställer konen på cirkeln på hennes röda cirkel .
han tar hennes blåa pil .
han tar hennes röda pil .
