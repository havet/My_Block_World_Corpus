
\data\
ngram 1= 35
ngram 2= 140
ngram 3= 294

\1-grams:
-3.33965	<s>	-2.10115
-1.65391	ta	-1.48495
-1.79558	det	-2.08189
-1.15924	röda	-2.17898
-1.51357	blocket	-2.36689
-0.894825	</s>
-1.43656	ställ	-1.70407
-1.35288	konen	-2.52859
-0.899529	på	-2.43933
-1.14237	den	-2.73997
-0.974162	cirkeln	-2.90862
-1.63208	han	-2.24736
-1.5876	tar	-1.47934
-2.17828	sitt	-1.38917
-1.57622	block	-2.30374
-1.64945	hon	-2.22981
-1.36193	ställer	-1.70659
-1.93311	sin	-1.76592
-1.31027	blåa	-1.96936
-1.6962	cirkel	-2.18256
-1.80817	en	-1.67117
-2.27895	blå	-1.40937
-2.12217	pil	-1.74819
-1.62365	jag	-2.25588
-2.27895	hennes	-1.18752
-1.9164	kon	-1.95904
-2.12217	ett	-1.5721
-2.64068	blått	-1.49831
-2.13553	pilen	-1.7344
-2.31846	hans	-1.24304
-2.1092	min	-1.46052
-2.41023	röd	-1.27107
-2.09661	mitt	-1.59843
-3.16356	rött	-0.845098
-2.09661	<unk>

\2-grams:
-0.765989	<s> ta	-1.28444
-0.546353	<s> ställ	-1.50356
-0.743876	<s> han	-2.10265
-0.761475	<s> hon	-2.0851
-0.735336	<s> jag	-2.11117
-0.571248	ta det	-1.5133
-0.783323	ta blocket	-1.30245
-0.730542	ta konen	-1.3536
-1.0309	ta den	-1.05257
-1.30438	ta en	-0.167658
-1.54598	ta hennes
-1.09364	ta ett	-1.00142
-1.54495	ta pilen	-0.876483
-1.41063	ta hans	-0.222085
-2.11379	ta min
-1.54461	ta mitt	-0.331399
-0.337052	det röda	-1.90451
-0.273683	det blåa	-1.96756
-0.977913	röda blocket	-1.60348
-0.991414	röda konen	-1.58969
-0.287086	röda cirkeln	-2.29146
-1.18406	röda block	-1.39936
-0.88062	röda cirkel	-1.70039
-1.34207	röda kon	-1.00041
-1.53905	röda pilen	-1.3536
-0.482505	blocket </s>
-0.175506	blocket på	-1.41891
-0.884073	ställ det	-1.42055
-0.773091	ställ blocket	-1.83072
-0.590165	ställ konen	-2.01215
-0.658065	ställ den	-1.6424
-1.03222	ställ en	-0.834443
-1.96315	ställ hennes	-0.700392
-1.76396	ställ ett	-0.331399
-1.37291	ställ pilen	-1.24446
-2.33844	ställ hans
-1.62867	ställ min	-0.700392
-1.76373	ställ mitt	-0.331399
-0.841715	konen </s>
-0.0686362	konen på	-1.74131
-0.386527	på den	-2.45244
-0.365749	på cirkeln	-2.47308
-1.16359	på sin	-1.67812
-1.46747	på en	-1.20099
-1.85248	på hennes	-1.00142
-2.06606	på hans	-0.553248
-1.51687	på min	-1.15269
-0.205219	den röda	-2.2145
-0.425997	den blåa	-1.99412
-0.147347	cirkeln </s>
-0.542427	cirkeln på	-1.64768
-0.463628	han tar	-0.725299
-0.186498	han ställer	-1.21891
-1.01685	tar det	-1.13972
-1.28369	tar blocket	-0.876483
-0.796872	tar konen	-1.3536
-1.09585	tar den	-1.05257
-0.97959	tar sitt	-1.00142
-1.37183	tar sin	-0.318995
-1.05923	tar en	-0.658352
-1.29077	tar hennes	-0.331399
-1.29013	tar ett	-0.632429
-1.47618	tar pilen	-0.456338
-1.2909	tar hans	-0.52351
-1.37315	tar min	-0.444329
-0.911104	tar mitt	-1.06837
-0.766506	sitt röda	-1.09833
-0.309026	sitt block	-1.24446
-0.556724	sitt blåa	-1.30245
-1.5917	sitt blått
-0.338171	block </s>
-0.269806	block på	-1.26192
-0.43375	hon tar	-0.764644
-0.203303	hon ställer	-1.12368
-1.2441	ställer det	-1.13972
-1.10538	ställer blocket	-1.57545
-0.675716	ställer konen	-2.00142
-0.732619	ställer den	-1.6424
-1.07949	ställer sitt	-0.862472
-1.44667	ställer sin	-0.94343
-1.02672	ställer en	-1.17751
-1.83969	ställer hennes	-0.331399
-1.1079	ställer ett	-0.92145
-1.60055	ställer pilen	-1.09833
-1.7045	ställer hans	-0.456338
-1.51731	ställer min	-0.876483
-1.13835	ställer mitt	-1.06837
-0.210791	sin röda	-1.58969
-0.501517	sin blåa	-1.30245
-1.26365	sin kon	-0.876483
-0.762717	blåa blocket	-1.66653
-0.676949	blåa konen	-1.75154
-0.483549	blåa cirkeln	-1.94343
-0.900651	blåa block	-1.5297
-1.15928	blåa cirkel	-1.03037
-1.75649	blåa pil	-0.456338
-1.25864	blåa kon	-1.17751
-1.89206	blåa pilen	-0.876483
-0.0542311	cirkel </s>
-0.9489	cirkel på	-0.553248
-0.83738	en cirkel	-1.39936
-0.489179	en blå	-1.26466
-0.721415	en pil	-1.21228
-1.0678	en kon	-0.876483
-0.629627	en röd	-1.12636
-0.584152	blå cirkel	-1.17751
-0.354723	blå pil	-0.854278
-0.584672	blå kon	-1.17751
-0.561305	pil </s>
-0.147476	pil på	-1.28397
-0.402932	jag tar	-1.0579
-0.222277	jag ställer	-1.19175
-0.350608	hennes röda	-0.745359
-0.768138	hennes block	-0.456338
-0.662613	hennes blåa	-0.553248
-1.10111	hennes cirkel	-0.700392
-1.48204	hennes pil
-0.644597	kon </s>
-0.11627	kon på	-1.18796
-0.167949	ett block	-1.44075
-0.617744	ett blått	-1.30245
-1.27092	ett rött	-0.700392
-0.0136334	blått block	-1.05257
-1.04621	pilen </s>
-0.0475309	pilen på	-0.942541
-0.721991	hans röda	-0.456338
-0.862549	hans block	-0.331399
-0.358019	hans blåa	-1.05257
-0.728474	hans cirkel	-0.456338
-0.348444	min röda	-1.27442
-0.575503	min blåa	-1.05257
-0.690029	min cirkel	-1.24446
-1.28094	min kon
-0.767712	röd cirkel	-0.876483
-0.633489	röd pil	-1.00142
-0.26337	röd kon	-1.3536
-0.588297	mitt röda	-1.3536
-0.393586	mitt block	-1.24446
-0.499819	mitt blåa	-1.44075
-0.0650307	rött block	-0.700392

\3-grams:
-0.551878	<s> ta det
-0.766828	<s> ta blocket
-0.714425	<s> ta konen
-1.02487	<s> ta den
-1.29664	<s> ta en
-1.54402	<s> ta hennes
-1.079	<s> ta ett
-1.54397	<s> ta pilen
-1.40306	<s> ta hans
-1.54395	<s> ta mitt
-0.873985	<s> ställ det
-0.762978	<s> ställ blocket
-0.579363	<s> ställ konen
-0.648763	<s> ställ den
-1.02345	<s> ställ en
-1.98244	<s> ställ hennes
-1.7721	<s> ställ ett
-1.36808	<s> ställ pilen
-1.63102	<s> ställ min
-1.77209	<s> ställ mitt
-0.461801	<s> han tar
-0.183987	<s> han ställer
-0.431738	<s> hon tar
-0.200726	<s> hon ställer
-0.400937	<s> jag tar
-0.21989	<s> jag ställer
-0.336942	ta det röda
-0.268043	ta det blåa
-0.308486	ta blocket </s>
-0.293837	ta blocket på
-0.26778	ta konen </s>
-0.33713	ta konen på
-0.246807	ta den röda
-0.363143	ta den blåa
-0.422036	ta en kon
-0.114713	ta ett block
-0.649368	ta ett blått
-0.00602532	ta pilen på
-0.178296	ta hans blåa
-0.166684	ta mitt blåa
-0.00486888	det röda blocket
-0.00388879	det blåa blocket
-0.363267	röda blocket </s>
-0.246666	röda blocket på
-1.05741	röda konen </s>
-0.0398496	röda konen på
-0.131788	röda cirkeln </s>
-0.582146	röda cirkeln på
-0.188179	röda block </s>
-0.454092	röda block på
-0.0667016	röda cirkel </s>
-0.846872	röda cirkel på
-0.0103123	röda kon på
-0.00199899	röda pilen på
-0.241868	blocket på den
-0.533373	blocket på cirkeln
-1.26508	blocket på sin
-1.51531	blocket på en
-1.52936	blocket på hans
-1.7178	blocket på min
-0.369511	ställ det röda
-0.242101	ställ det blåa
-0.00213734	ställ blocket på
-0.000617958	ställ konen på
-0.311112	ställ den röda
-0.291207	ställ den blåa
-0.450728	ställ en blå
-0.39661	ställ en pil
-0.682416	ställ en röd
-0.0508178	ställ hennes röda
-0.189638	ställ ett blått
-0.00257182	ställ pilen på
-0.310077	ställ min röda
-0.343608	ställ min blåa
-0.18437	ställ mitt röda
-0.373439	konen på den
-0.337295	konen på cirkeln
-1.18379	konen på sin
-1.46136	konen på en
-1.78735	konen på min
-0.16071	på den röda
-0.509629	på den blåa
-0.170169	på cirkeln </s>
-0.489217	på cirkeln på
-0.163274	på sin röda
-0.505971	på sin blåa
-0.288626	på en cirkel
-0.501393	på en blå
-0.819069	på en röd
-0.128064	på hennes röda
-0.68181	på hennes cirkel
-0.112082	på hans cirkel
-0.376903	på min röda
-0.765187	på min blåa
-0.395044	på min cirkel
-0.804788	den röda konen
-0.0985228	den röda cirkeln
-1.35595	den röda pilen
-0.42009	den blåa konen
-0.226821	den blåa cirkeln
-1.65414	den blåa pilen
-0.462696	cirkeln på den
-0.261179	cirkeln på cirkeln
-1.442	cirkeln på sin
-1.69195	cirkeln på en
-1.29827	cirkeln på min
-1.19478	han tar det
-1.25534	han tar blocket
-0.660235	han tar konen
-1.21576	han tar den
-0.745291	han tar sitt
-0.830063	han tar en
-1.07585	han tar ett
-1.0936	han tar pilen
-1.16209	han tar mitt
-1.23651	han ställer det
-1.1281	han ställer blocket
-0.691062	han ställer konen
-0.694412	han ställer den
-0.920089	han ställer sitt
-1.14341	han ställer sin
-0.975925	han ställer en
-1.12826	han ställer ett
-1.25119	han ställer pilen
-1.5428	han ställer mitt
-0.345187	tar det röda
-0.26137	tar det blåa
-0.507746	tar blocket </s>
-0.161821	tar blocket på
-0.186489	tar konen </s>
-0.457166	tar konen på
-0.632352	tar den röda
-0.115374	tar den blåa
-0.631083	tar sitt röda
-0.364145	tar sitt block
-0.484432	tar sitt blåa
-0.262486	tar sin kon
-0.47974	tar en blå
-0.554524	tar en kon
-0.506324	tar en röd
-0.46042	tar hennes block
-0.43383	tar hennes blåa
-0.0337475	tar ett block
-0.166365	tar pilen </s>
-0.489852	tar hans röda
-0.248018	tar hans blåa
-0.381118	tar min blåa
-0.469689	tar min kon
-0.553956	tar mitt röda
-0.439875	tar mitt block
-0.448925	tar mitt blåa
-0.0336329	sitt röda block
-0.673763	sitt block </s>
-0.103564	sitt block på
-0.019348	sitt blåa block
-0.36112	block på den
-0.512211	block på cirkeln
-0.799659	block på sin
-1.35831	block på en
-1.57518	block på hennes
-1.5608	block på min
-0.840574	hon tar det
-1.14311	hon tar konen
-0.84893	hon tar den
-0.760419	hon tar sitt
-0.969239	hon tar sin
-0.845225	hon tar en
-1.28599	hon tar min
-0.916731	hon tar mitt
-1.19842	hon ställer det
-1.31385	hon ställer blocket
-0.566022	hon ställer konen
-0.625446	hon ställer den
-0.883143	hon ställer sitt
-1.5385	hon ställer sin
-0.938205	hon ställer en
-1.18772	hon ställer ett
-1.49866	hon ställer mitt
-0.265544	ställer det röda
-0.340177	ställer det blåa
-0.00385492	ställer blocket på
-0.000632797	ställer konen på
-0.337285	ställer den röda
-0.2676	ställer den blåa
-0.908054	ställer sitt röda
-0.218276	ställer sitt block
-0.579762	ställer sitt blåa
-0.233154	ställer sin röda
-0.389859	ställer sin blåa
-0.410853	ställer en blå
-0.571462	ställer en pil
-0.485752	ställer en röd
-0.197119	ställer hennes blåa
-0.103392	ställer ett block
-0.693974	ställer ett blått
-0.00360517	ställer pilen på
-0.0949261	ställer hans blåa
-0.180591	ställer min röda
-0.5197	ställer min blåa
-0.865105	ställer mitt röda
-0.187825	ställer mitt block
-0.671955	ställer mitt blåa
-0.081323	sin röda cirkel
-0.82507	sin röda kon
-0.137549	sin blåa cirkel
-0.645979	sin blåa pil
-0.0470981	sin kon </s>
-0.270139	blåa blocket </s>
-0.334352	blåa blocket på
-1.21927	blåa konen </s>
-0.0270561	blåa konen på
-0.103401	blåa cirkeln </s>
-0.673957	blåa cirkeln på
-0.20175	blåa block </s>
-0.430075	blåa block på
-0.00478043	blåa cirkel </s>
-0.046086	blåa pil på
-0.634816	blåa kon </s>
-0.114856	blåa kon på
-0.00602532	blåa pilen på
-0.236097	cirkel på cirkeln
-0.578298	cirkel på hennes
-0.00203774	en cirkel </s>
-0.570621	en blå cirkel
-0.336822	en blå pil
-0.570648	en blå kon
-0.853809	en pil </s>
-0.0659251	en pil på
-0.200423	en kon </s>
-0.433484	en kon på
-0.756109	en röd cirkel
-0.61535	en röd pil
-0.237813	en röd kon
-0.0034011	blå cirkel </s>
-0.0178524	blå pil på
-0.00683183	blå kon på
-0.128923	pil på den
-0.868054	pil på cirkeln
-0.933046	pil på sin
-1.01657	jag tar det
-1.16749	jag tar blocket
-0.650219	jag tar konen
-1.33654	jag tar den
-0.932902	jag tar hennes
-1.36108	jag tar ett
-0.850484	jag tar hans
-1.36894	jag tar min
-0.70744	jag tar mitt
-1.34082	jag ställer det
-0.952656	jag ställer blocket
-0.733869	jag ställer konen
-0.871265	jag ställer den
-1.19292	jag ställer en
-1.36768	jag ställer hennes
-1.02064	jag ställer ett
-1.22654	jag ställer hans
-1.03481	jag ställer min
-0.797141	jag ställer mitt
-0.565598	hennes röda block
-0.233743	hennes röda cirkel
-0.0910684	hennes block </s>
-0.121808	hennes blåa block
-0.0102836	hennes cirkel </s>
-0.466391	kon på den
-0.28569	kon på cirkeln
-1.3518	kon på sin
-1.03506	kon på en
-0.38976	ett block </s>
-0.227488	ett block på
-0.000669704	ett blått block
-0.0122096	ett rött block
-0.481878	blått block </s>
-0.173945	blått block på
-0.675293	pilen på den
-0.146604	pilen på cirkeln
-1.21709	pilen på min
-0.171846	hans röda block
-0.126228	hans block </s>
-0.38586	hans blåa block
-0.287232	hans blåa kon
-0.161364	hans cirkel på
-0.34961	min röda cirkel
-0.293135	min röda kon
-0.529922	min blåa cirkel
-0.202558	min blåa kon
-0.0029134	min cirkel </s>
-0.00682912	röd cirkel </s>
-0.0325942	röd pil </s>
-0.00454244	röd kon på
-0.0183623	mitt röda block
-0.673763	mitt block </s>
-0.103564	mitt block på
-0.0139847	mitt blåa block
-0.0420302	rött block på
\end\
