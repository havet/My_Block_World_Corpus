ta det röda blocket .
ta blocket .
ställ konen på den röda cirkeln på cirkeln .
han tar sitt röda block .
hon ställer det röda blocket på sin blåa cirkel .
han ställer en blå pil på den röda cirkeln på en cirkel .
hon ställer det blåa blocket på den blåa cirkeln .
jag ställer hennes blåa kon på cirkeln på cirkeln .
han ställer sin blåa pil på den röda cirkeln .
hon ställer konen på cirkeln på cirkeln .
han tar ett blått block .
ställ den röda konen på den blåa cirkeln på cirkeln .
ställ det röda blocket på den blåa cirkeln .
ställ den blåa pilen på den blåa cirkeln .
ställ hennes röda kon på den blåa cirkeln på cirkeln .
ta hans block .
han ställer den röda konen på cirkeln på cirkeln .
han ställer konen på cirkeln på cirkeln .
jag ställer hans block på den blåa cirkeln på cirkeln .
jag tar det röda blocket .
jag tar konen på den röda cirkeln .
jag tar min kon på den röda cirkeln .
ställ konen på den röda cirkeln på hennes cirkel .
jag ställer en röd kon på cirkeln .
jag ställer min röda kon på cirkeln .
jag ställer min röda kon på min cirkel .
jag ställer konen på cirkeln på min cirkel .
han tar ett block .
jag ställer konen på den röda cirkeln på min röda cirkel .
hon ställer mitt blåa block på den blåa cirkeln .
hon tar min blåa kon .
han tar ett block på cirkeln .
hon tar pilen .
hon tar det röda blocket .
jag tar hans röda block .
han ställer konen på den röda cirkeln .
ställ den blåa konen på den röda cirkeln .
hon ställer den blåa konen på den blåa cirkeln .
han ställer den röda konen på den röda cirkeln .
han ställer sitt blåa block på sin röda cirkel .
jag ställer min blåa kon på den röda cirkeln .
jag ställer ett block på cirkeln på den röda cirkeln .
jag ställer mitt block på min cirkel .
jag ställer hennes block på min cirkel .
hon tar konen .
han tar en röd pil .
hon ställer sitt block på den röda cirkeln .
ställ pilen på den röda cirkeln på cirkeln .
hon ställer konen på sin röda cirkel på cirkeln .
ta konen på cirkeln .
jag ställer den blåa konen på den röda cirkeln på cirkeln .
hon ställer blocket på sin röda cirkel .
han ställer blocket på den blåa cirkeln .
hon tar det röda blocket på den blåa cirkeln .
han tar konen på sin röda cirkel .
jag ställer den blåa konen på den blåa cirkeln .
jag ställer det blåa blocket på den blåa cirkeln .
hon ställer konen på min röda cirkel på den röda cirkeln .
ställ det röda blocket på cirkeln på den blåa cirkeln .
jag tar hans blåa kon .
jag ställer blocket på den röda cirkeln .
jag tar mitt block .
jag ställer mitt block på den röda cirkeln .
ta konen på hans röda cirkel .
ställ hennes röda block på den röda cirkeln .
jag ställer blocket på den blåa cirkeln .
hon ställer blocket på cirkeln på sin blåa cirkel .
hon tar en röd pil .
jag ställer den röda pilen på hennes cirkel .
han ställer mitt röda block på en blå cirkel .
ställ en kon på den röda cirkeln på den röda cirkeln .
han ställer en pil på sin röda cirkel på cirkeln .
han tar sitt block på den röda cirkeln .
ta mitt blåa block .
ställ konen på den röda cirkeln på min cirkel .
han ställer sitt block på cirkeln på sin röda cirkel .
ställ konen på den blåa cirkeln .
han ställer konen på cirkeln på cirkeln .
han tar min röda kon på cirkeln .
hon ställer konen på cirkeln på den röda cirkeln .
ställ min blåa kon på cirkeln .
ställ konen på cirkeln .
han ställer konen på cirkeln .
hon ställer sitt blåa block på sin blåa cirkel .
hon tar sitt block .
hon tar mitt block .
ställ ett blått block på den röda cirkeln .
hon ställer pilen på cirkeln på den röda cirkeln .
han ställer den blåa konen på cirkeln .
han ställer en blå kon på en blå cirkel .
ställ blocket på den röda cirkeln .
han ställer den blåa konen på cirkeln på cirkeln .
han ställer den röda pilen på cirkeln .
hon ställer en blå pil på den blåa cirkeln .
ta pilen på cirkeln .
jag tar ett block .
jag tar mitt blåa block .
jag tar mitt röda block .
hon tar sitt blåa block .
jag ställer ett block på den blåa cirkeln på cirkeln .
jag ställer hans blåa kon på cirkeln .
han tar blocket på cirkeln .
hon tar sin kon .
hon ställer ett block på sin röda cirkel .
jag tar mitt röda block .
ställ min blåa kon på cirkeln .
han ställer sin blåa pil på sin röda cirkel .
hon tar sin kon .
hon tar det röda blocket .
han tar sitt blåa block .
jag tar hennes block .
jag ställer min röda kon på cirkeln .
hon ställer mitt block på cirkeln på den röda cirkeln .
ta ett block .
jag ställer konen på cirkeln på den röda cirkeln .
jag ställer den röda pilen på min cirkel .
hon ställer sitt röda block på sin röda cirkel .
ställ konen på cirkeln .
hon ställer ett rött block på en blå cirkel .
han ställer ett blått block på den röda cirkeln .
jag tar mitt blåa block .
jag tar konen .
han tar konen .
jag tar hennes blåa block .
ställ pilen på cirkeln på den röda cirkeln .
hon ställer den blåa konen på min blåa cirkel .
hon tar ett block på den röda cirkeln .
hon tar det blåa blocket .
jag ställer konen på cirkeln på cirkeln .
ta den röda konen på cirkeln .
han tar sitt röda block .
jag ställer hans blåa kon på den röda cirkeln .
jag ställer den blåa konen på cirkeln .
hon ställer den blåa konen på den röda cirkeln .
han ställer den blåa pilen på den blåa cirkeln .
ta hans blåa block .
ställ det röda blocket på den röda cirkeln .
jag tar den blåa konen på den röda cirkeln .
jag ställer mitt block på hennes röda cirkel .
hon ställer blocket på den röda cirkeln .
ta hans röda block .
ställ konen på den blåa cirkeln på cirkeln .
jag ställer en röd kon på cirkeln .
ställ en blå pil på den röda cirkeln på en cirkel .
jag ställer konen på den röda cirkeln på cirkeln .
jag ställer mitt blåa block på den blåa cirkeln .
han ställer en pil på den röda cirkeln på cirkeln .
ställ mitt blåa block på den röda cirkeln .
jag tar konen .
hon tar mitt blåa block .
hon tar den blåa konen .
han ställer den röda konen på en cirkel .
hon ställer konen på den röda cirkeln på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
jag ställer mitt röda block på den blåa cirkeln .
jag tar mitt blåa block .
ta ett block .
jag tar hennes blåa block .
jag ställer ett block på cirkeln på den blåa cirkeln .
hon ställer den röda konen på cirkeln på cirkeln .
ta den röda konen .
hon tar den blåa konen på den röda cirkeln .
han tar en blå pil .
ta blocket .
hon ställer konen på cirkeln på min röda cirkel .
hon ställer sin röda kon på den röda cirkeln .
hon tar en pil .
han tar en röd pil .
han tar pilen på cirkeln .
han ställer konen på cirkeln på min röda cirkel .
ställ mitt röda block på cirkeln .
hon ställer konen på den röda cirkeln på sin röda cirkel .
hon ställer den blåa konen på den röda cirkeln på cirkeln .
ta det blåa blocket .
hon tar min kon .
jag tar blocket på cirkeln .
jag tar hans block .
jag tar hans röda block .
ta min röda kon på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
ställ blocket på den blåa cirkeln på cirkeln .
ställ det blåa blocket på den röda cirkeln .
hon ställer det blåa blocket på sin blåa cirkel .
ta det röda blocket på den blåa cirkeln .
han ställer det blåa blocket på min blåa cirkel .
ta mitt röda block .
han tar den blåa konen på den röda cirkeln .
hon tar den röda konen .
ställ det blåa blocket på den blåa cirkeln .
han ställer sitt blått block på sin röda cirkel .
jag tar det blåa blocket .
ta det blåa blocket .
hon ställer den blåa konen på cirkeln .
han ställer den röda konen på den blåa cirkeln på cirkeln .
ta mitt blåa block .
ställ den blåa konen på cirkeln på cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta konen .
han ställer sin röda kon på cirkeln .
hon ställer konen på sin röda cirkel .
han ställer konen på sin röda cirkel på sin röda cirkel .
hon ställer konen på cirkeln på cirkeln .
hon tar konen på sin röda cirkel .
hon ställer sitt blåa block på sin röda cirkel .
han ställer konen på den röda cirkeln på cirkeln .
hon tar sin röda kon .
jag ställer ett block på den röda cirkeln .
han ställer mitt blåa block på sin blåa cirkel .
hon tar mitt block på cirkeln .
han ställer sitt block på cirkeln på den röda cirkeln .
hon ställer den blåa konen på sin röda cirkel .
ställ den röda konen på den röda cirkeln .
han tar en kon .
han ställer konen på sin blåa cirkel .
han ställer ett block på cirkeln på sin blåa cirkel .
han ställer den blåa konen på sin röda cirkel .
han ställer sitt blåa block på den blåa cirkeln .
han ställer blocket på sin blåa cirkel på cirkeln .
ställ en blå pil på cirkeln .
ta konen på den röda cirkeln .
hon tar sitt block .
jag tar konen .
jag tar min blåa kon på den blåa cirkeln .
hon ställer en röd kon på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
jag tar konen .
hon tar blocket på sin röda cirkel .
han ställer konen på cirkeln .
hon ställer sitt block på den blåa cirkeln .
han ställer en pil på den röda cirkeln .
hon tar sitt block på cirkeln .
jag ställer hans blåa block på den röda cirkeln .
hon ställer konen på cirkeln .
han ställer konen på cirkeln .
han tar sin blåa pil .
ta hennes röda block .
han ställer sitt block på sin röda cirkel .
han tar det blåa blocket .
han ställer blocket på cirkeln på cirkeln .
ta hennes block .
hon ställer det röda blocket på den blåa cirkeln .
han ställer den blåa konen på den blåa cirkeln .
jag ställer konen på den röda cirkeln på cirkeln .
han ställer ett block på den röda cirkeln .
jag tar den röda konen på cirkeln .
hon tar en kon .
jag tar det blåa blocket .
han tar det röda blocket .
ställ en röd kon på cirkeln .
ta blocket på hans cirkel .
jag tar hennes pil .
han ställer pilen på cirkeln på den röda cirkeln .
ta hans blåa kon .
hon ställer den blåa konen på sin röda cirkel .
jag ställer hennes blåa block på den blåa cirkeln .
han tar sitt block .
han ställer pilen på sin röda cirkel på cirkeln .
hon tar sitt röda block .
han tar hennes röda block .
han ställer konen på sin röda cirkel på cirkeln .
han tar pilen .
jag ställer mitt block på cirkeln på cirkeln .
han tar konen .
jag ställer min blåa kon på den blåa cirkeln .
ta blocket på cirkeln .
jag tar konen på cirkeln .
ställ pilen på cirkeln på den röda cirkeln .
hon ställer ett block på cirkeln på min blåa cirkel .
hon ställer en blå pil på sin blåa cirkel .
ta konen .
ställ en röd kon på cirkeln .
ställ mitt röda block på den blåa cirkeln .
jag ställer konen på cirkeln på den röda cirkeln .
han ställer den röda pilen på cirkeln på cirkeln .
ställ konen på cirkeln .
ställ blocket på cirkeln på cirkeln .
jag ställer konen på den röda cirkeln på den röda cirkeln .
ställ den röda konen på cirkeln .
jag tar hans blåa block .
han tar konen .
ställ konen på cirkeln på cirkeln .
ta det röda blocket .
jag tar mitt block på cirkeln .
han tar mitt röda block .
hon tar det blåa blocket .
ställ en pil på den röda cirkeln .
hon ställer en pil på den röda cirkeln på cirkeln .
hon ställer konen på cirkeln på cirkeln .
han ställer den blåa konen på den röda cirkeln .
han ställer sin röda kon på sin röda cirkel .
ställ blocket på den röda cirkeln .
han tar sitt blåa block .
hon tar mitt röda block .
han tar den blåa konen .
hon ställer den röda konen på cirkeln .
jag tar ett block .
ställ blocket på en röd cirkel .
jag tar konen .
hon ställer sitt block på den blåa cirkeln på cirkeln .
ta det blåa blocket .
jag ställer det röda blocket på den röda cirkeln .
han ställer blocket på min röda cirkel .
jag ställer ett block på hennes röda cirkel .
jag tar hans blåa block .
ställ blocket på den röda cirkeln .
jag ställer konen på cirkeln .
han tar en blå kon på den blåa cirkeln .
jag tar konen .
han ställer den blåa konen på den röda cirkeln på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
hon tar en kon .
ställ blocket på cirkeln på cirkeln .
hon ställer den blåa konen på den röda cirkeln på cirkeln .
han ställer ett blått block på sin röda cirkel .
han tar blocket .
han tar konen .
hon ställer konen på cirkeln .
hon tar sitt blåa block .
hon tar den blåa konen på sin blåa cirkel .
jag ställer blocket på den röda cirkeln .
jag tar blocket på den röda cirkeln .
hon ställer konen på cirkeln på sin röda cirkel .
jag ställer konen på den röda cirkeln på cirkeln .
jag ställer ett block på hans cirkel på hennes röda cirkel .
jag ställer min röda kon på den röda cirkeln .
ställ en pil på den röda cirkeln på cirkeln .
han ställer konen på en cirkel .
hon ställer den röda pilen på cirkeln .
jag tar hennes block .
jag tar mitt block .
han tar pilen .
hon ställer konen på cirkeln .
ställ blocket på cirkeln på den röda cirkeln .
han ställer det röda blocket på den blåa cirkeln .
ställ hans blåa kon på den blåa cirkeln .
jag ställer mitt block på den blåa cirkeln på cirkeln .
han ställer blocket på en röd cirkel .
ställ den röda pilen på cirkeln på cirkeln .
han ställer en blå pil på cirkeln .
jag ställer blocket på hans cirkel på hennes röda cirkel .
jag ställer den röda konen på den röda cirkeln .
jag ställer mitt block på cirkeln på cirkeln .
ta en kon på en cirkel .
han ställer det röda blocket på cirkeln .
jag ställer blocket på cirkeln på den röda cirkeln .
hon ställer sin röda kon på cirkeln .
jag tar konen på cirkeln .
jag ställer konen på den röda cirkeln på cirkeln .
hon ställer konen på en cirkel .
han ställer sitt block på cirkeln .
hon ställer ett block på sin blåa cirkel .
hon ställer konen på den röda cirkeln på den röda cirkeln .
hon ställer den röda konen på min röda cirkel .
ta ett blått block .
jag ställer det blåa blocket på den röda cirkeln .
hon ställer den röda konen på en cirkel .
han ställer en pil på den röda cirkeln på den röda cirkeln .
ställ konen på cirkeln på den röda cirkeln .
han ställer pilen på cirkeln på den röda cirkeln .
han tar mitt blåa block .
ställ min röda kon på den röda cirkeln .
jag ställer den röda konen på den blåa cirkeln på cirkeln .
han ställer pilen på cirkeln på min röda cirkel .
jag ställer en röd kon på cirkeln .
hon ställer sitt block på cirkeln .
ställ min röda kon på cirkeln .
hon ställer den blåa konen på cirkeln på cirkeln .
hon tar en blå kon på sin blåa cirkel .
han ställer det röda blocket på cirkeln på den blåa cirkeln .
hon ställer en blå kon på en blå cirkel .
ta hennes blåa block .
han ställer konen på cirkeln på den röda cirkeln .
han tar konen på cirkeln .
hon tar den blåa konen på den röda cirkeln .
ta ett block .
ställ konen på den röda cirkeln på cirkeln .
ta konen på cirkeln .
ta blocket .
ta ett block .
ställ en röd kon på cirkeln .
ställ blocket på den blåa cirkeln på cirkeln .
ställ den blåa konen på den blåa cirkeln .
ställ den blåa konen på den röda cirkeln .
ställ det blåa blocket på den röda cirkeln .
ställ det röda blocket på den röda cirkeln .
ställ den röda konen på den blåa cirkeln på cirkeln .
ta den blåa konen på den röda cirkeln .
ta den blåa konen på den blåa cirkeln .
ställ blocket på cirkeln på den röda cirkeln .
ta konen .
ta blocket .
ställ blocket på cirkeln på cirkeln .
ta det blåa blocket .
ta ett blått block .
ta konen på den röda cirkeln .
ställ blocket på den röda cirkeln .
ställ blocket på cirkeln på den röda cirkeln .
ta konen .
ställ den röda konen på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta blocket på cirkeln .
ta det röda blocket .
ta den röda konen på cirkeln .
ställ konen på den röda cirkeln på den röda cirkeln .
ställ blocket på den röda cirkeln .
ta det blåa blocket .
ställ blocket på den röda cirkeln .
ställ den blåa konen på den röda cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta konen .
ställ konen på den röda cirkeln på cirkeln .
ta det blåa blocket .
ställ konen på cirkeln på den röda cirkeln .
ställ konen på cirkeln på cirkeln .
ta blocket på den röda cirkeln .
ta blocket .
ställ den röda konen på den röda cirkeln .
ta det blåa blocket .
ta blocket .
ta det blåa blocket .
ställ den blåa konen på cirkeln .
ställ blocket på cirkeln på den blåa cirkeln .
ställ konen på den röda cirkeln på den röda cirkeln .
ta det röda blocket .
ställ den blåa konen på den blåa cirkeln .
ställ det röda blocket på den blåa cirkeln .
ställ konen på cirkeln .
ställ den blåa konen på cirkeln på cirkeln .
ställ konen på den röda cirkeln på cirkeln .
ställ det blåa blocket på den röda cirkeln .
ställ konen på den röda cirkeln på cirkeln .
ta konen .
ställ den blåa konen på cirkeln .
ta konen .
ställ den blåa konen på den röda cirkeln på cirkeln .
ställ den röda konen på den röda cirkeln .
ställ blocket på den blåa cirkeln .
ta konen på cirkeln .
ställ konen på cirkeln på cirkeln .
ställ blocket på den röda cirkeln .
ta blocket på cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta det röda blocket .
ta konen .
ställ konen på cirkeln .
ta den röda konen .
ställ konen på cirkeln på den röda cirkeln .
ställ den röda konen på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
ta det röda blocket på den blåa cirkeln .
ta det röda blocket .
ta blocket .
ställ det röda blocket på den blåa cirkeln .
ställ blocket på cirkeln på cirkeln .
ställ konen på cirkeln på den röda cirkeln .
ställ det röda blocket på cirkeln .
ställ konen på cirkeln .
ställ blocket på den blåa cirkeln på cirkeln .
ställ konen på den röda cirkeln .
ta det röda blocket .
ställ det röda blocket på cirkeln på den blåa cirkeln .
ställ konen på den röda cirkeln på cirkeln .
ställ den blåa konen på den blåa cirkeln .
ställ blocket på cirkeln .
ställ konen på cirkeln .
ta det blåa blocket .
ställ den röda konen på cirkeln på cirkeln .
ställ blocket på den röda cirkeln .
ställ den blåa konen på den röda cirkeln .
ställ den röda konen på cirkeln .
ställ den blåa konen på den röda cirkeln på cirkeln .
ta den blåa konen .
ställ det röda blocket på den blåa cirkeln .
ställ det blåa blocket på den röda cirkeln .
ställ konen på den blåa cirkeln .
ta det blåa blocket .
ställ en pil på den röda cirkeln på cirkeln .
ta pilen på cirkeln .
ta ett block .
jag ställer en röd kon på cirkeln .
hon ställer en röd kon på cirkeln .
jag ställer mitt block på den blåa cirkeln på cirkeln .
hon ställer en blå pil på den blåa cirkeln .
han ställer sin blåa pil på den röda cirkeln .
han ställer ett blått block på den röda cirkeln .
hon ställer sitt röda block på den röda cirkeln .
ställ den röda konen på den blåa cirkeln på cirkeln .
ta den blåa konen på den röda cirkeln .
ta en blå kon på den blåa cirkeln .
han ställer sitt block på cirkeln på den röda cirkeln .
han tar konen .
jag tar blocket .
jag ställer mitt block på cirkeln på cirkeln .
jag tar det blåa blocket .
ta konen på den röda cirkeln .
jag ställer blocket på hennes röda cirkel .
jag ställer blocket på hans cirkel på hennes röda cirkel .
hon tar sin kon .
jag ställer den röda pilen på min cirkel .
ställ konen på cirkeln på den röda cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta blocket på cirkeln .
ta det röda blocket .
ta den röda konen på cirkeln .
ställ en pil på den röda cirkeln på den röda cirkeln .
ställ blocket på en röd cirkel .
ta det blåa blocket .
ställ blocket på den röda cirkeln .
ställ den blåa konen på den röda cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta konen .
ställ pilen på den röda cirkeln på cirkeln .
ta det blåa blocket .
ställ pilen på cirkeln på den röda cirkeln .
ställ konen på cirkeln på cirkeln .
ta blocket på den röda cirkeln .
ta ett block .
ställ den röda konen på den röda cirkeln .
ta det blåa blocket .
ta blocket .
ta det blåa blocket .
ställ den blåa konen på cirkeln .
ställ blocket på cirkeln på den blåa cirkeln .
ställ konen på den röda cirkeln på den röda cirkeln .
ta det röda blocket .
ställ en blå kon på en blå cirkel .
ställ ett rött block på en blå cirkel .
ställ konen på en cirkel .
ställ den blåa konen på cirkeln på cirkeln .
ställ en pil på den röda cirkeln på cirkeln .
ställ ett blått block på den röda cirkeln .
ställ konen på den röda cirkeln på cirkeln .
ta konen .
ställ en blå pil på cirkeln .
ta en kon .
ställ en blå pil på den röda cirkeln på en cirkel .
ställ den röda konen på den röda cirkeln .
ställ blocket på den blåa cirkeln .
ta konen på cirkeln .
ställ konen på cirkeln på cirkeln .
ställ blocket på den röda cirkeln .
ta blocket på cirkeln .
ställ det blåa blocket på den blåa cirkeln .
ta det röda blocket .
ta pilen på cirkeln .
ställ konen på cirkeln .
ta en röd pil .
ställ den röda pilen på cirkeln .
ställ pilen på cirkeln på den röda cirkeln .
ställ pilen på cirkeln på den röda cirkeln .
ställ den blåa pilen på den blåa cirkeln .
ställ den röda pilen på cirkeln på cirkeln .
ställ en pil på den röda cirkeln .
ställ den röda konen på en cirkel .
ta en pil .
